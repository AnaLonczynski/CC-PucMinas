/*
 Guia_0205.v
 680668 - Ana Clara Lonczynski
*/
module Guia_0205;
// define data
  reg [7:0] a1 = 8'b101_110, b1 = 8'b1000_101, C1 = 8'b101_101, d1 = 8'b10111_01, e1 = 8'b1101011; // binary
  reg [7:0] a2 = 8'b10_011, b2 = 8'b10_010, c2 = 8'b10_101, d2 = 8'b11_011, e2 = 8'b1101; // binary
  reg [7:0] c1;
 initial
 begin : main
   $display ( "\nGuia_0205 - Tests" );
 c1 = a1+a2;
 $display ( "\na.) 101,11(2) + 10,011(2) = %8b", c1 );
 c1 = b1-b2;
 $display ( "\nb.) 1000,101(2) - 10,01(2) = %8b", c1 );
 c1 = C1*c2;
 $display ( "\nc.) 101,101(2) * 10,101(2) = %8b", c1 );
 c1 = d1/d2;
 $display ( "\nd.) 10111,01(2) / 11,011(2) = %8b", c1 );
 c1 = e1%e2;
   $display ( "\ne.) 1101011(2) % 1101(2) = %8b", c1 );
 end // main
endmodule // Guia_0205

/*SAIDA:
Guia_0205 - Tests

a.) 101,11(2) + 10,011(2) = 01000001

b.) 1000,101(2) - 10,01(2) = 00110011

c.) 101,101(2) * 10,101(2) = 10110001

d.) 10111,01(2) / 11,011(2) = 00000011

e.) 1101011(2) % 1101(2) = 00000011
*/